interface iterate_page_i;
endinterface
