module iterate_page ();
endmodule
